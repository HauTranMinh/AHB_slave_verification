package AHB_slave_pkg;

	`include "C:/Users/LENOVO/Desktop/AHB/AHB_slave/AHB_slave_transaction.sv";
	`include "C:/Users/LENOVO/Desktop/AHB/AHB_slave/AHB_types.sv";
	`include "C:/Users/LENOVO/Desktop/AHB/AHB_slave/AHB_slave_sequencer.sv";
	`include "C:/Users/LENOVO/Desktop/AHB/AHB_slave/AHB_slave_sequence_read.sv";
	`include "C:/Users/LENOVO/Desktop/AHB/AHB_slave/AHB_slave_sequence_write.sv";
	`include "C:/Users/LENOVO/Desktop/AHB/AHB_slave/AHB_slave_driver.sv";
	`include "C:/Users/LENOVO/Desktop/AHB/AHB_slave/AHB_slave_monitor.sv";
	`include "C:/Users/LENOVO/Desktop/AHB/AHB_slave/AHB_slave_agent.sv";



endpackage