 class AHB_types extends uvm_object;
 	
 endclass : AHB_types